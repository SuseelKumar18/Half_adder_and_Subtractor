// Half Subtractor in Verilog 
module half_subtractor ( 
    input  wire a, b,         // Inputs 
    output wire diff, borrow  // Outputs 
); 
 
    // Logic equations 
    assign diff   = a ^ b;     // XOR for difference 
    assign borrow = ~a & b;    // Borrow when a < b 
 
endmodule 